
/*
This module is a latch-based control system for addressing within the
accumulator table. Since The addressing for each column of the accumulator table
is the same in successive clock cycles (column M writes to address A in clock
cycle N, and column M+1 writes to address A in clock cycle N+1), it is only
necessary to control the addressing of the first column. The addressing of the
first column is passed along the pipeline, where a column receives the address
from the column to its left in the following clock cycle.
*/

module accumTableWr_control (clk,
                             reset,
                             wr_en_in,
                             data_mem_calc_done,
                             sub_row,
                             submat_m,
                             submat_n,
                             wr_en_out,
                             wr_addr_out);

    parameter MAX_OUT_ROWS = 128; // output number of rows in 
    parameter MAX_OUT_COLS = 128;
    parameter SYS_ARR_ROWS = 16;
    parameter SYS_ARR_COLS = 16;
    
    localparam NUM_ACCUM_ROWS = MAX_OUT_ROWS * (MAX_OUT_COLS/SYS_ARR_COLS);
    localparam ADDR_WIDTH = $clog2(NUM_ACCUM_ROWS);
    localparam NUM_SUBMATS_M = MAX_OUT_ROWS/SYS_ARR_ROWS; // not sure if this will do ceiling like I want
    localparam NUM_SUBMATS_N = MAX_OUT_COLS/SYS_ARR_COLS; // not sure if this will do ceiling like I want

    input clk;
    input reset;
    input wr_en_in;
    input data_mem_calc_done;
    input [$clog2(SYS_ARR_ROWS)-1:0] sub_row;
    input [$clog2(NUM_SUBMATS_M)-1:0] submat_m; // sub-matrix row number (sub-matrix position in the overall matrix)
    input [$clog2(NUM_SUBMATS_N)-1:0] submat_n; // sub-matrix col number (sub-matrix position in the overall matrix)
    output wire [SYS_ARR_COLS-1:0] wr_en_out; // LSB is first column
    output wire [ADDR_WIDTH*SYS_ARR_COLS-1:0] wr_addr_out; // LSBs are first column

    wire [ADDR_WIDTH-1:0] addr_0;
    reg [SYS_ARR_COLS-2:0] wr_en_out_partial, wr_en_out_partial_c;
    reg [ADDR_WIDTH*(SYS_ARR_COLS-1)-1:0] wr_addr_out_partial, wr_addr_out_partial_c;
    reg [$clog2(SYS_ARR_ROWS)-1:0] count_c, count;

    accumTableAddr_control accumTableAddr_control (
        .sub_row (sub_row),
        .submat_m(submat_m),
        .submat_n(submat_n),
        .addr    (addr_0)
    );

    assign wr_en_out = (data_mem_calc_done == 1) ? {wr_en_out_partial, wr_en_in} : {SYS_ARR_COLS{8'hx}};
    assign wr_addr_out = (data_mem_calc_done == 1) ? {wr_addr_out_partial, addr_0} : {SYS_ARR_COLS * ADDR_WIDTH {8'hx}};
    assign sub_row = count;
    
    always @(clk, reset, wr_en_in, sub_row, submat_m, submat_n) begin
        
        if((wr_en_in) && (count_c < 16)) begin
            count_c = count + 4'b0001;
        end
        else begin
            count_c = 4'b0000;
        end
        
        wr_en_out_partial_c[0] = wr_en_in;
        wr_addr_out_partial_c[ADDR_WIDTH-1:0] = addr_0;
        
        wr_en_out_partial_c[SYS_ARR_COLS-1:1] = wr_en_out_partial[SYS_ARR_COLS-2:0];
        wr_addr_out_partial_c[ADDR_WIDTH*(SYS_ARR_COLS-1)-1:ADDR_WIDTH] = wr_addr_out_partial[ADDR_WIDTH*(SYS_ARR_COLS-2)-1:0];
        
       
        if (reset) begin
                    wr_en_out_partial_c = {SYS_ARR_COLS-1{1'b0}};
                    count_c = {($clog2(SYS_ARR_ROWS) + 1){1'b0}};
                    count = {($clog2(SYS_ARR_ROWS) + 1){1'b0}};
        end // if (reset)
    end // always @(clk, reset, wr_en_in, sub_row, submat_m, submat_n) 

    always @(posedge clk) begin
        wr_en_out_partial <= wr_en_out_partial_c;
        wr_addr_out_partial <= wr_addr_out_partial_c;
        count <= count_c;
    end // always @(posedge clk)

endmodule
